// NOR gates.
//f(A, B, C, D)= ∑m(0,1,2,5,8,9,10)

module q2(a, b, c, d, f);
    input a, b, c, d;
    output f;
    wire g0, g1, g2, g3, g4, g5, g6, g7;


